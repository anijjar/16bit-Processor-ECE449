
-- 2:1 MuX
X <= A when S = '1' else B;